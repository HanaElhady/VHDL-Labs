library ieee;
use ieee.std_logic_1164.all;

entity assign_4 is 
	port(
	x,y : in std_logic_vector(3 downto 0);	
	cin : in std_logic;
	sum : out std_logic_vector(3 downto 0);
	cout : out std_logic
	);									 
end assign_4 ;




